library verilog;
use verilog.vl_types.all;
entity testBench_lcdController is
end testBench_lcdController;
