module LCDcontrollerTop
(

);


endmodule
